LIBRARY 	ieee;
USE		ieee.std_logic_1164.all, ieee.numeric_std.all;

ENTITY de10liteg IS
	PORT(	
		CLOCK_50	: IN	std_logic;
		KEY		: IN 	std_logic_vector( 1 DOWNTO 0 );
		SW			: IN 	std_logic_vector( 9 DOWNTO 0 );
		GPIO_24	: IN	std_logic;	--RX
		GPIO_25	: OUT std_logic;	--TX
		LEDR		: OUT	std_logic_vector( 9 DOWNTO 0 )
	);
END de10liteg;

ARCHITECTURE Structural OF de10liteg IS	
	
	component gumnut_with_mem IS
		generic( 
			IMem_file_name	: string 	:= "gasm_text.dat";
			DMem_file_name : string 	:= "gasm_data.dat";
         debug 			: boolean	:= false 
		);
		port( 
			clk_i 			: in 	std_logic;
         rst_i 			: in 	std_logic;
         -- I/O port bus
         port_cyc_o 		: out	std_logic;
         port_stb_o 		: out std_logic;
         port_we_o 		: out std_logic;
         port_ack_i 		: in 	std_logic;
         port_adr_o 		: out unsigned(7 downto 0);
         port_dat_o 		: out std_logic_vector(7 downto 0);
         port_dat_i 		: in 	std_logic_vector(7 downto 0);
         -- Interrupts
         int_req 			: in std_logic;
         int_ack 			: out std_logic
		);
	end component gumnut_with_mem;
	
	COMPONENT uart IS
		GENERIC(
			clk_freq  	: integer    := 50_000_000;  	--frequency of system clock in Hertz
			baud_rate 	: integer    := 115_200;     	--data link baud rate in bits/second
			os_rate   	: integer    := 16;          	--oversampling rate to find center of receive bits (in samples per baud period)
			d_width   	: integer    := 8;           	--data bus width
			parity    	: integer    := 0;           	--0 for no parity, 1 for parity
			parity_eo	: std_logic  := '0'				--'0' for even, '1' for odd parity
		);        
		PORT(
			clk      	: IN  std_logic;                             --system clock
			reset_n		: IN  std_logic;                             --ascynchronous reset
			tx_ena   	: IN  std_logic;                             --initiate transmission
			tx_data  	: IN  std_logic_vector(d_width-1 DOWNTO 0);  --data to transmit
			rx       	: IN  std_logic;                             --receive pin
			rx_busy  	: OUT std_logic;                             --data reception in progress, LEDR(9)
			rx_error 	: OUT std_logic;                             --start, parity, or stop bit error detected
			rx_data  	: OUT std_logic_vector(d_width-1 DOWNTO 0);  --data received
			tx_busy  	: OUT std_logic;                             --transmission in progress, LEDR(8)
			tx       	: OUT	std_logic										--transmit pin
		);                            
	END COMPONENT;

	COMPONENT debounce IS
		PORT(	
			Clock			: IN		std_logic;
			button		: IN		std_logic;
			debounced	: BUFFER	std_logic
		);
	END COMPONENT;
	
	SIGNAL clk_i, rst_i				: std_logic; 
	SIGNAL port_cyc_o, port_stb_o	: std_logic;
	SIGNAL port_we_o, port_ack_i	: std_logic;
	SIGNAL int_req, int_ack			: std_logic;
	SIGNAL port_adr_o					: unsigned(7 DOWNTO 0);
	SIGNAL port_dat_o, port_dat_i	: std_logic_vector(7 DOWNTO 0);
	
	SIGNAL tx_ena_de10						: std_logic	:= '1';
	SIGNAL tx_data_de10, rx_data_de10	: std_logic_vector(7 DOWNTO 0);
	SIGNAL rx_busy_de10, rx_error_de10	: std_logic;
	SIGNAL tx_busy_de10						: std_logic;
	
	SIGNAL key1_db			: std_logic;
	
BEGIN
	rst_i	<= not KEY( 0 );
	LEDR 	<= ( OTHERS => '0' );
	
	gumnut		: gumnut_with_mem 
						PORT MAP(
								CLOCK_50, 
								rst_i, 
								port_cyc_o, 
								port_stb_o, 
								port_we_o, 
								'1', 
								port_adr_o,
								port_dat_o, 
								port_dat_i,
								int_req, 
								int_ack
						);

	uart_de10	: uart 		
						PORT MAP( 
								CLOCK_50, 
								KEY(0), 
								tx_ena_de10, 
								tx_data_de10, 
								GPIO_24, 
								rx_busy_de10, 
								rx_error_de10, 
								rx_data_de10, 
								tx_busy_de10, 
								GPIO_25 
						);
	
	button_de10	: debounce	
						PORT MAP( 
								CLOCK_50, 
								KEY(1), 
								key1_db 
						);	
	
	-- Output => TX_DATA -> data memory address: 0x00
	PROCESS( CLOCK_50, rst_i )
		BEGIN
			IF rst_i = '1' THEN
				tx_data_de10 <= ( OTHERS => '0' );
			ELSIF rising_edge( CLOCK_50 ) THEN	
				IF port_adr_o 	= "00000000"	and	-- address port 
					port_cyc_o 	= '1' 			and	-- control signals for I/O
					port_stb_o 	= '1' 			and 
					port_we_o  	= '1'					-- 'write' operation 			
				THEN	
					tx_data_de10 <= port_dat_o;
				END IF;
			END IF;
	END PROCESS;
	
	-- Output => TX_START -> data memory address: 0x01
	PROCESS( CLOCK_50, rst_i )
		BEGIN
			IF rst_i = '1' THEN
				tx_ena_de10 <= '1';
			ELSIF rising_edge( CLOCK_50 ) THEN	
				IF port_adr_o 	= "00000001"	and	-- address port 
					port_cyc_o 	= '1' 			and	-- control signals for I/O
					port_stb_o 	= '1' 			and 
					port_we_o  	= '1'					-- 'write' operation 			
				THEN	
					tx_ena_de10 <= port_dat_o(0);
				END IF;
			END IF;
	END PROCESS;
	
	-- Input <= KEY1 -> data memory address: 0x02
	PROCESS( CLOCK_50, rst_i )
		BEGIN
			IF rst_i = '1' THEN
				port_dat_i <= ( OTHERS => '0' );
			ELSIF rising_edge( CLOCK_50 ) THEN 
				IF port_adr_o		= "00000011"	and	-- address port 
					port_cyc_o 		= '1' 			and	-- control signals for I/O
					port_stb_o 		= '1' 			and 
					port_we_o  		= '0'						-- 'read' operation
				THEN	
					port_dat_i <= "0000000" & key1_db;
				END IF;	
			END IF;
	END PROCESS;
		
END Structural;